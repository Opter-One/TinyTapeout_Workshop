/*
 * Copyright (c) 2024 Uri Shaked
 * SPDX-License-Identifier: Apache-2.0
 */

`default_nettype none

module tt_um_Opter_One_VGA_direction(
  input  wire [7:0] ui_in,    // Dedicated inputs
  output wire [7:0] uo_out,   // Dedicated outputs
  input  wire [7:0] uio_in,   // IOs: Input path
  output wire [7:0] uio_out,  // IOs: Output path
  output wire [7:0] uio_oe,   // IOs: Enable path (active high: 0=input, 1=output)
  input  wire       ena,      // always 1 when the design is powered, so you can ignore it
  input  wire       clk,      // clock
  input  wire       rst_n     // reset_n - low to reset
);

  // VGA signals
  wire hsync;
  wire vsync;
  wire [1:0] R;
  wire [1:0] G;
  wire [1:0] B;
  wire video_active;
  wire [9:0] pix_x;
  wire [9:0] pix_y;
  wire sound;

  // TinyVGA PMOD
  assign uo_out = {hsync, B[0], G[0], R[0], vsync, B[1], G[1], R[1]};

  // Unused outputs assigned to 0.
  assign uio_out = 0;
  assign uio_oe  = 0;

  // Suppress unused signals warning
  wire _unused_ok = &{ena, ui_in, uio_in};

  reg [9:0] counter_x;
  reg [9:0] counter_y;
  reg [9:0] direction_y = 1;
  reg [9:0] direction_x = 1;

  hvsync_generator hvsync_gen(
    .clk(clk),
    .reset(~rst_n),
    .hsync(hsync),
    .vsync(vsync),
    .display_on(video_active),
    .hpos(pix_x),
    .vpos(pix_y)
  );
  
  wire [9:0] moving_x = pix_x + counter_x;
  wire [9:0] moving_y = pix_y + counter_y;

  assign R = video_active ? {moving_x[5], moving_y[5]} : 2'b00;
  assign G = video_active ? {moving_x[6], moving_y[6]} : 2'b00;
  assign B = video_active ? {moving_x[7], moving_y[7]} : 2'b00;
  
  always @(posedge vsync, negedge rst_n) begin
    if (~rst_n) begin
      counter_x <= 0;
      counter_y <= 0;
    end else begin

      if(counter_y == 256) begin
        direction_y <= -1;
      end if(counter_y == 0) begin
        direction_y <= 1;
      end

      if(counter_x == 512) begin
        direction_x <= -1;
      end if(counter_x == 0) begin
        direction_x <= 1;
      end
      
      counter_x <= counter_x + direction_x;
      counter_y <= counter_y + 2*direction_y;
      
    end
  end
  
endmodule
